`define RTMLAMP_OHWR_REGS_SIZE 1024
`define ADDR_RTMLAMP_OHWR_REGS_STA 'h0
`define RTMLAMP_OHWR_REGS_STA_RESERVED_OFFSET 0
`define RTMLAMP_OHWR_REGS_STA_RESERVED 'hffffffff
`define ADDR_RTMLAMP_OHWR_REGS_CTL 'h4
`define RTMLAMP_OHWR_REGS_CTL_RESERVED_OFFSET 0
`define RTMLAMP_OHWR_REGS_CTL_RESERVED 'hffffffff
`define ADDR_RTMLAMP_OHWR_REGS_CH 'h200
`define RTMLAMP_OHWR_REGS_CH_SIZE 512
`define ADDR_RTMLAMP_OHWR_REGS_CH_0 'h200
`define RTMLAMP_OHWR_REGS_CH_0_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_0_STA 'h200
`define RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_0_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_0_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_0_CTL 'h204
`define RTMLAMP_OHWR_REGS_CH_0_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_0_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_0_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_0_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_0_PI_KP 'h208
`define RTMLAMP_OHWR_REGS_CH_0_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_0_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_0_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_0_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_0_PI_TI 'h20c
`define RTMLAMP_OHWR_REGS_CH_0_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_0_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_0_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_0_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_0_PI_SP 'h210
`define RTMLAMP_OHWR_REGS_CH_0_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_0_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_0_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_0_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_0_DAC 'h214
`define RTMLAMP_OHWR_REGS_CH_0_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_0_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_0_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_0_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_0_LIM 'h218
`define RTMLAMP_OHWR_REGS_CH_0_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_0_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_0_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_0_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_0_CNT 'h21c
`define RTMLAMP_OHWR_REGS_CH_0_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_0_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_0_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_0_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_1 'h220
`define RTMLAMP_OHWR_REGS_CH_1_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_1_STA 'h220
`define RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_1_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_1_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_1_CTL 'h224
`define RTMLAMP_OHWR_REGS_CH_1_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_1_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_1_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_1_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_1_PI_KP 'h228
`define RTMLAMP_OHWR_REGS_CH_1_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_1_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_1_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_1_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_1_PI_TI 'h22c
`define RTMLAMP_OHWR_REGS_CH_1_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_1_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_1_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_1_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_1_PI_SP 'h230
`define RTMLAMP_OHWR_REGS_CH_1_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_1_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_1_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_1_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_1_DAC 'h234
`define RTMLAMP_OHWR_REGS_CH_1_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_1_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_1_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_1_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_1_LIM 'h238
`define RTMLAMP_OHWR_REGS_CH_1_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_1_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_1_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_1_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_1_CNT 'h23c
`define RTMLAMP_OHWR_REGS_CH_1_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_1_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_1_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_1_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_2 'h240
`define RTMLAMP_OHWR_REGS_CH_2_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_2_STA 'h240
`define RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_2_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_2_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_2_CTL 'h244
`define RTMLAMP_OHWR_REGS_CH_2_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_2_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_2_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_2_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_2_PI_KP 'h248
`define RTMLAMP_OHWR_REGS_CH_2_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_2_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_2_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_2_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_2_PI_TI 'h24c
`define RTMLAMP_OHWR_REGS_CH_2_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_2_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_2_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_2_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_2_PI_SP 'h250
`define RTMLAMP_OHWR_REGS_CH_2_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_2_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_2_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_2_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_2_DAC 'h254
`define RTMLAMP_OHWR_REGS_CH_2_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_2_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_2_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_2_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_2_LIM 'h258
`define RTMLAMP_OHWR_REGS_CH_2_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_2_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_2_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_2_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_2_CNT 'h25c
`define RTMLAMP_OHWR_REGS_CH_2_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_2_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_2_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_2_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_3 'h260
`define RTMLAMP_OHWR_REGS_CH_3_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_3_STA 'h260
`define RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_3_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_3_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_3_CTL 'h264
`define RTMLAMP_OHWR_REGS_CH_3_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_3_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_3_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_3_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_3_PI_KP 'h268
`define RTMLAMP_OHWR_REGS_CH_3_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_3_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_3_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_3_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_3_PI_TI 'h26c
`define RTMLAMP_OHWR_REGS_CH_3_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_3_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_3_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_3_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_3_PI_SP 'h270
`define RTMLAMP_OHWR_REGS_CH_3_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_3_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_3_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_3_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_3_DAC 'h274
`define RTMLAMP_OHWR_REGS_CH_3_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_3_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_3_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_3_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_3_LIM 'h278
`define RTMLAMP_OHWR_REGS_CH_3_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_3_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_3_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_3_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_3_CNT 'h27c
`define RTMLAMP_OHWR_REGS_CH_3_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_3_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_3_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_3_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_4 'h280
`define RTMLAMP_OHWR_REGS_CH_4_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_4_STA 'h280
`define RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_4_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_4_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_4_CTL 'h284
`define RTMLAMP_OHWR_REGS_CH_4_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_4_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_4_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_4_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_4_PI_KP 'h288
`define RTMLAMP_OHWR_REGS_CH_4_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_4_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_4_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_4_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_4_PI_TI 'h28c
`define RTMLAMP_OHWR_REGS_CH_4_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_4_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_4_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_4_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_4_PI_SP 'h290
`define RTMLAMP_OHWR_REGS_CH_4_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_4_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_4_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_4_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_4_DAC 'h294
`define RTMLAMP_OHWR_REGS_CH_4_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_4_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_4_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_4_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_4_LIM 'h298
`define RTMLAMP_OHWR_REGS_CH_4_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_4_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_4_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_4_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_4_CNT 'h29c
`define RTMLAMP_OHWR_REGS_CH_4_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_4_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_4_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_4_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_5 'h2a0
`define RTMLAMP_OHWR_REGS_CH_5_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_5_STA 'h2a0
`define RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_5_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_5_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_5_CTL 'h2a4
`define RTMLAMP_OHWR_REGS_CH_5_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_5_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_5_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_5_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_5_PI_KP 'h2a8
`define RTMLAMP_OHWR_REGS_CH_5_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_5_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_5_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_5_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_5_PI_TI 'h2ac
`define RTMLAMP_OHWR_REGS_CH_5_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_5_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_5_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_5_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_5_PI_SP 'h2b0
`define RTMLAMP_OHWR_REGS_CH_5_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_5_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_5_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_5_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_5_DAC 'h2b4
`define RTMLAMP_OHWR_REGS_CH_5_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_5_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_5_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_5_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_5_LIM 'h2b8
`define RTMLAMP_OHWR_REGS_CH_5_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_5_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_5_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_5_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_5_CNT 'h2bc
`define RTMLAMP_OHWR_REGS_CH_5_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_5_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_5_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_5_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_6 'h2c0
`define RTMLAMP_OHWR_REGS_CH_6_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_6_STA 'h2c0
`define RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_6_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_6_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_6_CTL 'h2c4
`define RTMLAMP_OHWR_REGS_CH_6_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_6_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_6_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_6_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_6_PI_KP 'h2c8
`define RTMLAMP_OHWR_REGS_CH_6_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_6_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_6_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_6_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_6_PI_TI 'h2cc
`define RTMLAMP_OHWR_REGS_CH_6_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_6_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_6_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_6_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_6_PI_SP 'h2d0
`define RTMLAMP_OHWR_REGS_CH_6_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_6_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_6_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_6_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_6_DAC 'h2d4
`define RTMLAMP_OHWR_REGS_CH_6_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_6_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_6_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_6_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_6_LIM 'h2d8
`define RTMLAMP_OHWR_REGS_CH_6_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_6_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_6_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_6_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_6_CNT 'h2dc
`define RTMLAMP_OHWR_REGS_CH_6_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_6_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_6_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_6_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_7 'h2e0
`define RTMLAMP_OHWR_REGS_CH_7_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_7_STA 'h2e0
`define RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_7_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_7_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_7_CTL 'h2e4
`define RTMLAMP_OHWR_REGS_CH_7_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_7_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_7_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_7_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_7_PI_KP 'h2e8
`define RTMLAMP_OHWR_REGS_CH_7_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_7_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_7_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_7_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_7_PI_TI 'h2ec
`define RTMLAMP_OHWR_REGS_CH_7_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_7_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_7_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_7_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_7_PI_SP 'h2f0
`define RTMLAMP_OHWR_REGS_CH_7_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_7_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_7_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_7_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_7_DAC 'h2f4
`define RTMLAMP_OHWR_REGS_CH_7_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_7_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_7_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_7_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_7_LIM 'h2f8
`define RTMLAMP_OHWR_REGS_CH_7_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_7_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_7_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_7_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_7_CNT 'h2fc
`define RTMLAMP_OHWR_REGS_CH_7_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_7_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_7_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_7_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_8 'h300
`define RTMLAMP_OHWR_REGS_CH_8_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_8_STA 'h300
`define RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_8_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_8_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_8_CTL 'h304
`define RTMLAMP_OHWR_REGS_CH_8_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_8_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_8_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_8_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_8_PI_KP 'h308
`define RTMLAMP_OHWR_REGS_CH_8_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_8_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_8_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_8_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_8_PI_TI 'h30c
`define RTMLAMP_OHWR_REGS_CH_8_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_8_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_8_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_8_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_8_PI_SP 'h310
`define RTMLAMP_OHWR_REGS_CH_8_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_8_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_8_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_8_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_8_DAC 'h314
`define RTMLAMP_OHWR_REGS_CH_8_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_8_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_8_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_8_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_8_LIM 'h318
`define RTMLAMP_OHWR_REGS_CH_8_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_8_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_8_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_8_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_8_CNT 'h31c
`define RTMLAMP_OHWR_REGS_CH_8_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_8_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_8_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_8_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_9 'h320
`define RTMLAMP_OHWR_REGS_CH_9_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_9_STA 'h320
`define RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_9_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_9_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_9_CTL 'h324
`define RTMLAMP_OHWR_REGS_CH_9_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_9_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_9_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_9_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_9_PI_KP 'h328
`define RTMLAMP_OHWR_REGS_CH_9_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_9_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_9_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_9_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_9_PI_TI 'h32c
`define RTMLAMP_OHWR_REGS_CH_9_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_9_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_9_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_9_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_9_PI_SP 'h330
`define RTMLAMP_OHWR_REGS_CH_9_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_9_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_9_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_9_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_9_DAC 'h334
`define RTMLAMP_OHWR_REGS_CH_9_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_9_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_9_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_9_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_9_LIM 'h338
`define RTMLAMP_OHWR_REGS_CH_9_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_9_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_9_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_9_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_9_CNT 'h33c
`define RTMLAMP_OHWR_REGS_CH_9_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_9_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_9_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_9_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_10 'h340
`define RTMLAMP_OHWR_REGS_CH_10_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_10_STA 'h340
`define RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_10_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_10_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_10_CTL 'h344
`define RTMLAMP_OHWR_REGS_CH_10_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_10_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_10_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_10_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_10_PI_KP 'h348
`define RTMLAMP_OHWR_REGS_CH_10_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_10_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_10_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_10_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_10_PI_TI 'h34c
`define RTMLAMP_OHWR_REGS_CH_10_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_10_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_10_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_10_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_10_PI_SP 'h350
`define RTMLAMP_OHWR_REGS_CH_10_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_10_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_10_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_10_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_10_DAC 'h354
`define RTMLAMP_OHWR_REGS_CH_10_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_10_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_10_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_10_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_10_LIM 'h358
`define RTMLAMP_OHWR_REGS_CH_10_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_10_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_10_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_10_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_10_CNT 'h35c
`define RTMLAMP_OHWR_REGS_CH_10_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_10_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_10_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_10_CNT_RESERVED 'hffc00000
`define ADDR_RTMLAMP_OHWR_REGS_CH_11 'h360
`define RTMLAMP_OHWR_REGS_CH_11_SIZE 32
`define ADDR_RTMLAMP_OHWR_REGS_CH_11_STA 'h360
`define RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_L_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_L 'h1
`define RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_L_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_L 'h2
`define RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_R_OFFSET 2
`define RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_R 'h4
`define RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_R_OFFSET 3
`define RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_R 'h8
`define RTMLAMP_OHWR_REGS_CH_11_STA_RESERVED_OFFSET 4
`define RTMLAMP_OHWR_REGS_CH_11_STA_RESERVED 'hfffffff0
`define ADDR_RTMLAMP_OHWR_REGS_CH_11_CTL 'h364
`define RTMLAMP_OHWR_REGS_CH_11_CTL_AMP_EN_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_11_CTL_AMP_EN 'h1
`define RTMLAMP_OHWR_REGS_CH_11_CTL_MODE_OFFSET 1
`define RTMLAMP_OHWR_REGS_CH_11_CTL_MODE 'h1e
`define ADDR_RTMLAMP_OHWR_REGS_CH_11_PI_KP 'h368
`define RTMLAMP_OHWR_REGS_CH_11_PI_KP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_11_PI_KP_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_11_PI_KP_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_11_PI_KP_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_11_PI_TI 'h36c
`define RTMLAMP_OHWR_REGS_CH_11_PI_TI_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_11_PI_TI_DATA 'h3ffffff
`define RTMLAMP_OHWR_REGS_CH_11_PI_TI_RESERVED_OFFSET 26
`define RTMLAMP_OHWR_REGS_CH_11_PI_TI_RESERVED 'hfc000000
`define ADDR_RTMLAMP_OHWR_REGS_CH_11_PI_SP 'h370
`define RTMLAMP_OHWR_REGS_CH_11_PI_SP_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_11_PI_SP_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_11_PI_SP_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_11_PI_SP_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_11_DAC 'h374
`define RTMLAMP_OHWR_REGS_CH_11_DAC_DATA_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_11_DAC_DATA 'hffff
`define RTMLAMP_OHWR_REGS_CH_11_DAC_RESERVED_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_11_DAC_RESERVED 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_11_LIM 'h378
`define RTMLAMP_OHWR_REGS_CH_11_LIM_LIM_A_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_11_LIM_LIM_A 'hffff
`define RTMLAMP_OHWR_REGS_CH_11_LIM_LIM_B_OFFSET 16
`define RTMLAMP_OHWR_REGS_CH_11_LIM_LIM_B 'hffff0000
`define ADDR_RTMLAMP_OHWR_REGS_CH_11_CNT 'h37c
`define RTMLAMP_OHWR_REGS_CH_11_CNT_CNT_OFFSET 0
`define RTMLAMP_OHWR_REGS_CH_11_CNT_CNT 'h3fffff
`define RTMLAMP_OHWR_REGS_CH_11_CNT_RESERVED_OFFSET 22
`define RTMLAMP_OHWR_REGS_CH_11_CNT_RESERVED 'hffc00000
