package rtmlamp_ohwr_regs_consts_pkg is
  constant c_RTMLAMP_OHWR_REGS_SIZE : Natural := 552;
  constant c_RTMLAMP_OHWR_REGS_STA_ADDR : Natural := 16#0#;
  constant c_RTMLAMP_OHWR_REGS_STA_RESERVED_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CTL_ADDR : Natural := 16#4#;
  constant c_RTMLAMP_OHWR_REGS_CTL_DAC_DATA_FROM_WB_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CTL_RESERVED_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_0_STA_ADDR : Natural := 16#100#;
  constant c_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_0_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_0_CTL_ADDR : Natural := 16#104#;
  constant c_RTMLAMP_OHWR_REGS_CH_0_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_0_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_0_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_0_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_0_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_0_PI_KP_ADDR : Natural := 16#108#;
  constant c_RTMLAMP_OHWR_REGS_CH_0_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_0_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_0_PI_TI_ADDR : Natural := 16#10c#;
  constant c_RTMLAMP_OHWR_REGS_CH_0_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_0_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_0_PI_SP_ADDR : Natural := 16#110#;
  constant c_RTMLAMP_OHWR_REGS_CH_0_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_0_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_0_DAC_ADDR : Natural := 16#114#;
  constant c_RTMLAMP_OHWR_REGS_CH_0_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_0_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_0_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_1_STA_ADDR : Natural := 16#118#;
  constant c_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_1_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_1_CTL_ADDR : Natural := 16#11c#;
  constant c_RTMLAMP_OHWR_REGS_CH_1_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_1_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_1_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_1_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_1_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_1_PI_KP_ADDR : Natural := 16#120#;
  constant c_RTMLAMP_OHWR_REGS_CH_1_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_1_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_1_PI_TI_ADDR : Natural := 16#124#;
  constant c_RTMLAMP_OHWR_REGS_CH_1_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_1_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_1_PI_SP_ADDR : Natural := 16#128#;
  constant c_RTMLAMP_OHWR_REGS_CH_1_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_1_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_1_DAC_ADDR : Natural := 16#12c#;
  constant c_RTMLAMP_OHWR_REGS_CH_1_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_1_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_1_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_2_STA_ADDR : Natural := 16#130#;
  constant c_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_2_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_2_CTL_ADDR : Natural := 16#134#;
  constant c_RTMLAMP_OHWR_REGS_CH_2_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_2_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_2_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_2_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_2_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_2_PI_KP_ADDR : Natural := 16#138#;
  constant c_RTMLAMP_OHWR_REGS_CH_2_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_2_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_2_PI_TI_ADDR : Natural := 16#13c#;
  constant c_RTMLAMP_OHWR_REGS_CH_2_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_2_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_2_PI_SP_ADDR : Natural := 16#140#;
  constant c_RTMLAMP_OHWR_REGS_CH_2_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_2_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_2_DAC_ADDR : Natural := 16#144#;
  constant c_RTMLAMP_OHWR_REGS_CH_2_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_2_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_2_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_3_STA_ADDR : Natural := 16#148#;
  constant c_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_3_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_3_CTL_ADDR : Natural := 16#14c#;
  constant c_RTMLAMP_OHWR_REGS_CH_3_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_3_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_3_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_3_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_3_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_3_PI_KP_ADDR : Natural := 16#150#;
  constant c_RTMLAMP_OHWR_REGS_CH_3_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_3_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_3_PI_TI_ADDR : Natural := 16#154#;
  constant c_RTMLAMP_OHWR_REGS_CH_3_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_3_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_3_PI_SP_ADDR : Natural := 16#158#;
  constant c_RTMLAMP_OHWR_REGS_CH_3_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_3_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_3_DAC_ADDR : Natural := 16#15c#;
  constant c_RTMLAMP_OHWR_REGS_CH_3_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_3_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_3_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_4_STA_ADDR : Natural := 16#160#;
  constant c_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_4_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_4_CTL_ADDR : Natural := 16#164#;
  constant c_RTMLAMP_OHWR_REGS_CH_4_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_4_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_4_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_4_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_4_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_4_PI_KP_ADDR : Natural := 16#168#;
  constant c_RTMLAMP_OHWR_REGS_CH_4_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_4_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_4_PI_TI_ADDR : Natural := 16#16c#;
  constant c_RTMLAMP_OHWR_REGS_CH_4_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_4_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_4_PI_SP_ADDR : Natural := 16#170#;
  constant c_RTMLAMP_OHWR_REGS_CH_4_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_4_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_4_DAC_ADDR : Natural := 16#174#;
  constant c_RTMLAMP_OHWR_REGS_CH_4_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_4_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_4_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_5_STA_ADDR : Natural := 16#178#;
  constant c_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_5_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_5_CTL_ADDR : Natural := 16#17c#;
  constant c_RTMLAMP_OHWR_REGS_CH_5_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_5_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_5_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_5_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_5_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_5_PI_KP_ADDR : Natural := 16#180#;
  constant c_RTMLAMP_OHWR_REGS_CH_5_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_5_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_5_PI_TI_ADDR : Natural := 16#184#;
  constant c_RTMLAMP_OHWR_REGS_CH_5_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_5_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_5_PI_SP_ADDR : Natural := 16#188#;
  constant c_RTMLAMP_OHWR_REGS_CH_5_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_5_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_5_DAC_ADDR : Natural := 16#18c#;
  constant c_RTMLAMP_OHWR_REGS_CH_5_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_5_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_5_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_6_STA_ADDR : Natural := 16#190#;
  constant c_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_6_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_6_CTL_ADDR : Natural := 16#194#;
  constant c_RTMLAMP_OHWR_REGS_CH_6_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_6_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_6_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_6_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_6_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_6_PI_KP_ADDR : Natural := 16#198#;
  constant c_RTMLAMP_OHWR_REGS_CH_6_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_6_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_6_PI_TI_ADDR : Natural := 16#19c#;
  constant c_RTMLAMP_OHWR_REGS_CH_6_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_6_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_6_PI_SP_ADDR : Natural := 16#1a0#;
  constant c_RTMLAMP_OHWR_REGS_CH_6_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_6_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_6_DAC_ADDR : Natural := 16#1a4#;
  constant c_RTMLAMP_OHWR_REGS_CH_6_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_6_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_6_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_7_STA_ADDR : Natural := 16#1a8#;
  constant c_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_7_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_7_CTL_ADDR : Natural := 16#1ac#;
  constant c_RTMLAMP_OHWR_REGS_CH_7_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_7_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_7_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_7_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_7_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_7_PI_KP_ADDR : Natural := 16#1b0#;
  constant c_RTMLAMP_OHWR_REGS_CH_7_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_7_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_7_PI_TI_ADDR : Natural := 16#1b4#;
  constant c_RTMLAMP_OHWR_REGS_CH_7_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_7_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_7_PI_SP_ADDR : Natural := 16#1b8#;
  constant c_RTMLAMP_OHWR_REGS_CH_7_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_7_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_7_DAC_ADDR : Natural := 16#1bc#;
  constant c_RTMLAMP_OHWR_REGS_CH_7_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_7_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_7_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_8_STA_ADDR : Natural := 16#1c0#;
  constant c_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_8_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_8_CTL_ADDR : Natural := 16#1c4#;
  constant c_RTMLAMP_OHWR_REGS_CH_8_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_8_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_8_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_8_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_8_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_8_PI_KP_ADDR : Natural := 16#1c8#;
  constant c_RTMLAMP_OHWR_REGS_CH_8_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_8_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_8_PI_TI_ADDR : Natural := 16#1cc#;
  constant c_RTMLAMP_OHWR_REGS_CH_8_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_8_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_8_PI_SP_ADDR : Natural := 16#1d0#;
  constant c_RTMLAMP_OHWR_REGS_CH_8_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_8_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_8_DAC_ADDR : Natural := 16#1d4#;
  constant c_RTMLAMP_OHWR_REGS_CH_8_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_8_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_8_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_9_STA_ADDR : Natural := 16#1d8#;
  constant c_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_9_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_9_CTL_ADDR : Natural := 16#1dc#;
  constant c_RTMLAMP_OHWR_REGS_CH_9_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_9_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_9_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_9_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_9_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_9_PI_KP_ADDR : Natural := 16#1e0#;
  constant c_RTMLAMP_OHWR_REGS_CH_9_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_9_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_9_PI_TI_ADDR : Natural := 16#1e4#;
  constant c_RTMLAMP_OHWR_REGS_CH_9_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_9_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_9_PI_SP_ADDR : Natural := 16#1e8#;
  constant c_RTMLAMP_OHWR_REGS_CH_9_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_9_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_9_DAC_ADDR : Natural := 16#1ec#;
  constant c_RTMLAMP_OHWR_REGS_CH_9_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_9_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_9_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_10_STA_ADDR : Natural := 16#1f0#;
  constant c_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_10_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_10_CTL_ADDR : Natural := 16#1f4#;
  constant c_RTMLAMP_OHWR_REGS_CH_10_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_10_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_10_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_10_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_10_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_10_PI_KP_ADDR : Natural := 16#1f8#;
  constant c_RTMLAMP_OHWR_REGS_CH_10_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_10_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_10_PI_TI_ADDR : Natural := 16#1fc#;
  constant c_RTMLAMP_OHWR_REGS_CH_10_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_10_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_10_PI_SP_ADDR : Natural := 16#200#;
  constant c_RTMLAMP_OHWR_REGS_CH_10_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_10_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_10_DAC_ADDR : Natural := 16#204#;
  constant c_RTMLAMP_OHWR_REGS_CH_10_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_10_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_10_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_CH_11_STA_ADDR : Natural := 16#208#;
  constant c_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_L_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_L_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_R_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_R_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_11_STA_RESERVED_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_11_CTL_ADDR : Natural := 16#20c#;
  constant c_RTMLAMP_OHWR_REGS_CH_11_CTL_AMP_EN_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_11_CTL_PI_OL_TRIANG_ENABLE_OFFSET : Natural := 1;
  constant c_RTMLAMP_OHWR_REGS_CH_11_CTL_PI_OL_SQUARE_ENABLE_OFFSET : Natural := 2;
  constant c_RTMLAMP_OHWR_REGS_CH_11_CTL_PI_SP_SQUARE_ENABLE_OFFSET : Natural := 3;
  constant c_RTMLAMP_OHWR_REGS_CH_11_CTL_PI_ENABLE_OFFSET : Natural := 4;
  constant c_RTMLAMP_OHWR_REGS_CH_11_PI_KP_ADDR : Natural := 16#210#;
  constant c_RTMLAMP_OHWR_REGS_CH_11_PI_KP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_11_PI_KP_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_11_PI_TI_ADDR : Natural := 16#214#;
  constant c_RTMLAMP_OHWR_REGS_CH_11_PI_TI_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_11_PI_TI_RESERVED_OFFSET : Natural := 26;
  constant c_RTMLAMP_OHWR_REGS_CH_11_PI_SP_ADDR : Natural := 16#218#;
  constant c_RTMLAMP_OHWR_REGS_CH_11_PI_SP_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_11_PI_SP_RESERVED_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_11_DAC_ADDR : Natural := 16#21c#;
  constant c_RTMLAMP_OHWR_REGS_CH_11_DAC_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_CH_11_DAC_WR_OFFSET : Natural := 16;
  constant c_RTMLAMP_OHWR_REGS_CH_11_DAC_RESERVED_OFFSET : Natural := 17;
  constant c_RTMLAMP_OHWR_REGS_PI_OL_DAC_CNT_MAX_ADDR : Natural := 16#220#;
  constant c_RTMLAMP_OHWR_REGS_PI_OL_DAC_CNT_MAX_DATA_OFFSET : Natural := 0;
  constant c_RTMLAMP_OHWR_REGS_PI_OL_DAC_CNT_MAX_RESERVED_OFFSET : Natural := 22;
  constant c_RTMLAMP_OHWR_REGS_PI_SP_LIM_INF_ADDR : Natural := 16#224#;
  constant c_RTMLAMP_OHWR_REGS_PI_SP_LIM_INF_DATA_OFFSET : Natural := 0;
end package rtmlamp_ohwr_regs_consts_pkg;
