`define WB_RTMLAMP_OHWR_REGS_SIZE 128
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH 'h0
`define WB_RTMLAMP_OHWR_REGS_CH_SIZE 128
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_0 'h0
`define WB_RTMLAMP_OHWR_REGS_CH_0_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_0_STA 'h0
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_0_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_0_CTL 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_0_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_0_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_0_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_0_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_1 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_1_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_1_STA 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_1_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_1_CTL 'hc
`define WB_RTMLAMP_OHWR_REGS_CH_1_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_1_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_1_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_1_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_2 'h10
`define WB_RTMLAMP_OHWR_REGS_CH_2_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_2_STA 'h10
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_2_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_2_CTL 'h14
`define WB_RTMLAMP_OHWR_REGS_CH_2_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_2_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_2_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_2_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_3 'h18
`define WB_RTMLAMP_OHWR_REGS_CH_3_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_3_STA 'h18
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_3_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_3_CTL 'h1c
`define WB_RTMLAMP_OHWR_REGS_CH_3_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_3_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_3_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_3_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_4 'h20
`define WB_RTMLAMP_OHWR_REGS_CH_4_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_4_STA 'h20
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_4_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_4_CTL 'h24
`define WB_RTMLAMP_OHWR_REGS_CH_4_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_4_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_4_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_4_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_5 'h28
`define WB_RTMLAMP_OHWR_REGS_CH_5_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_5_STA 'h28
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_5_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_5_CTL 'h2c
`define WB_RTMLAMP_OHWR_REGS_CH_5_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_5_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_5_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_5_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_6 'h30
`define WB_RTMLAMP_OHWR_REGS_CH_6_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_6_STA 'h30
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_6_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_6_CTL 'h34
`define WB_RTMLAMP_OHWR_REGS_CH_6_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_6_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_6_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_6_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_7 'h38
`define WB_RTMLAMP_OHWR_REGS_CH_7_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_7_STA 'h38
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_7_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_7_CTL 'h3c
`define WB_RTMLAMP_OHWR_REGS_CH_7_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_7_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_7_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_7_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_8 'h40
`define WB_RTMLAMP_OHWR_REGS_CH_8_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_8_STA 'h40
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_8_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_8_CTL 'h44
`define WB_RTMLAMP_OHWR_REGS_CH_8_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_8_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_8_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_8_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_9 'h48
`define WB_RTMLAMP_OHWR_REGS_CH_9_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_9_STA 'h48
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_9_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_9_CTL 'h4c
`define WB_RTMLAMP_OHWR_REGS_CH_9_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_9_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_9_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_9_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_10 'h50
`define WB_RTMLAMP_OHWR_REGS_CH_10_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_10_STA 'h50
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_10_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_10_CTL 'h54
`define WB_RTMLAMP_OHWR_REGS_CH_10_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_10_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_10_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_10_CTL_RESERVED 'hfffffffe
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_11 'h58
`define WB_RTMLAMP_OHWR_REGS_CH_11_SIZE 8
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_11_STA 'h58
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_L_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_L 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_L_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_L 'h2
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_R_OFFSET 2
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_IFLAG_R 'h4
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_R_OFFSET 3
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_AMP_TFLAG_R 'h8
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_RESERVED_OFFSET 4
`define WB_RTMLAMP_OHWR_REGS_CH_11_STA_RESERVED 'hfffffff0
`define ADDR_WB_RTMLAMP_OHWR_REGS_CH_11_CTL 'h5c
`define WB_RTMLAMP_OHWR_REGS_CH_11_CTL_AMP_EN_OFFSET 0
`define WB_RTMLAMP_OHWR_REGS_CH_11_CTL_AMP_EN 'h1
`define WB_RTMLAMP_OHWR_REGS_CH_11_CTL_RESERVED_OFFSET 1
`define WB_RTMLAMP_OHWR_REGS_CH_11_CTL_RESERVED 'hfffffffe
